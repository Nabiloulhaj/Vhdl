library ieee;
use ieee.std_logic_1164.all;

entity BaudClkGenerator_tb is
end entity;


architecture rtl of BaudClkGenerator_tb is

	component BaudClkGenerator is
	generic 
	(
		 NUMBER_OF_CLOCKS    : integer := 10;
		 SYS_CLK_FREQ        : integer := 50000000;
		 BAUD_RATE           : integer := 115200
	);
	port
	(
		 Clk : in std_logic; -- 50MHz
		 Rst : in std_logic;
		 Start   : in std_logic;
		 BaudClk : out std_logic;
		 Ready   : out std_logic
	);
	end component;
	
	signal Clks 		: std_logic := '0';
	signal Rsts 		: std_logic;
	signal Starts   	: std_logic;
	signal BaudClks 	: std_logic;
	signal Readys   	: std_logic;

begin
	
	-- clks <= not clk after 10ns;
	
	clkgen:process
	begin
		clks <= '0';
		wait for 10ns;
		clks <= '1';
		wait for 10ns;
	end process;
	
	UUT: BaudClkGenerator 
	generic map(NUMBER_OF_CLOCKS =>10,SYS_CLK_FREQ =>50000000,BAUD_RATE =>115200)
	port map(Clk => clks ,Rst => rsts , start => starts , Baudclk => baudclks , Ready => readys);

	main:process
	begin
		rsts <= '1'; 
		starts <= '0';
		wait for 50ns;
		rsts <= '0';
		
		wait until rising_edge(clks);
		starts <= '1';
		wait until rising_edge(clks);
		starts <= '0';
		
		
		wait; -- stop process for repeating itself
	
	end process;

end rtl;